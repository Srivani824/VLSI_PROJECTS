package router_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"

`include "src_xtn.sv"
`include "src_config.sv"
`include "dst_config.sv"
`include "env_config.sv"
`include "src_drv.sv"
`include "src_mon.sv"
`include "src_seqr.sv"
`include "src_agt.sv"
`include "src_agt_top.sv"
`include "src_seqs.sv"

`include "dst_xtn.sv"
`include "dst_mon.sv"
`include "dst_seqr.sv"
`include "dst_seqs.sv"
`include "dst_drv.sv"
`include "dst_agt.sv"
`include "dst_agt_top.sv"

`include "v_seqr.sv"
`include "v_seqs.sv"
`include "scoreboard.sv"

`include "env.sv"

`include "test.sv"

endpackage
